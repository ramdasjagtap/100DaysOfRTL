`timescale 1ns / 1ps

//printing "HELLO WORLD"  in system verilog by using class.
class Day22;

  function void hello_world();
   $display("Hello World! \n");
  endfunction
endclass